module cpu
import rv32i_types::*;
(
    input   logic           clk,
    input   logic           rst,

    output  logic   [31:0]  imem_addr,
    output  logic   [3:0]   imem_rmask,
    input   logic   [31:0]  imem_rdata,
    input   logic           imem_resp,

    output  logic   [31:0]  dmem_addr,
    output  logic   [3:0]   dmem_rmask,
    output  logic   [3:0]   dmem_wmask,
    input   logic   [31:0]  dmem_rdata,
    output  logic   [31:0]  dmem_wdata,
    input   logic           dmem_resp
);

    if_id_stage_reg_t   curr_if_id_stage_reg, next_if_id_stage_reg;
    id_ex_stage_reg_t   curr_id_ex_stage_reg, next_id_ex_stage_reg;
    ex_mem_stage_reg_t  curr_ex_mem_stage_reg, next_ex_mem_stage_reg;
    mem_wb_stage_reg_t  curr_mem_wb_stage_reg, next_mem_wb_stage_reg;
    logic               stall;
    logic [4:0]         wb_rd_s;
    logic [31:0]        wb_rd_v;
    logic               wb_regf_we;
    id_rs1_forward_sel_t         id_rs1_forward_sel;
    id_rs2_forward_sel_t         id_rs2_forward_sel;
    ex_rs1_forward_sel_t         ex_rs1_forward_sel;
    ex_rs2_forward_sel_t         ex_rs2_forward_sel;
    logic  [4:0]    id_rs1_s;
    logic  [4:0]    id_rs2_s;
    logic  need_flush;
    logic  [31:0]  target_pc;

    Forwarding forwarding(
        .id_rs1_s(id_rs1_s),
        .id_rs2_s(id_rs2_s),
        .id_ex_stage_reg(curr_id_ex_stage_reg),
        .ex_mem_stage_reg(curr_ex_mem_stage_reg),
        .mem_wb_stage_reg(curr_mem_wb_stage_reg),
        .stall(stall),
        .id_rs1_forward_sel(id_rs1_forward_sel),
        .id_rs2_forward_sel(id_rs2_forward_sel),
        .ex_rs1_forward_sel(ex_rs1_forward_sel),
        .ex_rs2_forward_sel(ex_rs2_forward_sel)
    );

    IF_Stage if_stage(
        .clk(clk),
        .rst(rst),
        .imem_addr(imem_addr),
        .imem_rmask(imem_rmask),
        .not_stall(~stall),
        .if_id_stage_reg(next_if_id_stage_reg),
        .need_flush(need_flush),
        .target_pc(target_pc)
    );

    always_ff @ (posedge clk ) begin 
        if (rst) begin 
            curr_if_id_stage_reg <= '0;
        end else if (~stall) begin 
            curr_if_id_stage_reg <= next_if_id_stage_reg;
        end 
    end 

    ID_Stage id_stage(
        .clk(clk),
        .rst(rst),
        .if_id_stage_reg(curr_if_id_stage_reg),
        .id_ex_stage_reg(next_id_ex_stage_reg),
        .imem_resp(imem_resp),
        .imem_rdata(imem_rdata),
        .wb_rd_s(wb_rd_s),
        .wb_rd_v(wb_rd_v),
        .wb_regf_we(wb_regf_we),
        .stall(stall),
        .id_rs1_s(id_rs1_s),
        .id_rs2_s(id_rs2_s),
        .id_rs1_forward_sel(id_rs1_forward_sel),
        .id_rs2_forward_sel(id_rs2_forward_sel),
        .need_flush(need_flush)
    );

    always_ff @ (posedge clk ) begin 
        if (rst) begin 
            curr_id_ex_stage_reg <= '0;
        end else begin 
            curr_id_ex_stage_reg <= next_id_ex_stage_reg;
        end 
    end

    EX_Stage ex_stage(
        .id_ex_stage_reg(curr_id_ex_stage_reg),
        .ex_mem_stage_reg(next_ex_mem_stage_reg),
        .ex_mem_stage_reg_curr(curr_ex_mem_stage_reg),
        .wb_rd_v(wb_rd_v),
        .ex_rs1_forward_sel(ex_rs1_forward_sel),
        .ex_rs2_forward_sel(ex_rs2_forward_sel),
        .need_flush(need_flush),
        .target_pc(target_pc)
    );

    always_ff @ (posedge clk ) begin 
        if (rst) begin 
            curr_ex_mem_stage_reg <= '0;
        end else begin 
            curr_ex_mem_stage_reg <= next_ex_mem_stage_reg;
        end 
    end

    MEM_Stage mem_stage(
        .dmem_addr(dmem_addr),
        .dmem_rmask(dmem_rmask),
        .dmem_wmask(dmem_wmask),
        .dmem_wdata(dmem_wdata),
        .ex_mem_stage_reg(curr_ex_mem_stage_reg),
        .mem_wb_stage_reg(next_mem_wb_stage_reg)
    );

    always_ff @ (posedge clk ) begin 
        if (rst) begin 
            curr_mem_wb_stage_reg <= '0;
        end else begin 
            curr_mem_wb_stage_reg <= next_mem_wb_stage_reg;
        end 
    end

    WB_Stage wb_stage(
        .mem_wb_stage_reg(curr_mem_wb_stage_reg),
        .dmem_resp(dmem_resp),
        .dmem_rdata(dmem_rdata),
        .wb_rd_s(wb_rd_s),
        .wb_rd_v(wb_rd_v),
        .wb_regf_we(wb_regf_we)
    );


endmodule : cpu
