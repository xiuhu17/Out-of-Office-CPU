package cache_types;


endpackage