// [way 3][way 2][way 1][way 0]
module HITMISS(
    input logic [23:0] dirty_tag_0,
    input logic [23:0] dirty_tag_1,
    input logic [23:0] dirty_tag_2,
    input logic [23:0] dirty_tag_3,
    input logic valid_0,
    input logic valid_1,
    input logic valid_2,
    input logic valid_3,
    input logic [23:0] curr_tag,
    output logic [3:0] way_mask,
    output logic hit
);


endmodule