module top(
    input   logic           clk,
    input   logic           rst,
    output  logic           ack
);

            logic           req;
            logic   [3:0]   req_key;

    a a(.*);
    b b(.*);

endmodule
