// module Forwarding(

// );


// endmodule : Forwarding