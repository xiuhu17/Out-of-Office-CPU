module PLRU(
    input logic clk,
    input logic rst,
    input logic hit,
    input logic ufp_Resp,
    input logic [3:0] curr_set,
    output logic [1:0] curr_way_replace
);



endmodule