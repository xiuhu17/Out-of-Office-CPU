module lfsr #(
  parameter bit [15:0] SEED_VALUE = 'hECEB
) (
  input               clk,
  input               rst,
  input               en,
  output logic        rand_bit,
  output logic [15:0] shift_reg
);

  // TODO: Fill this out!

endmodule : lfsr
