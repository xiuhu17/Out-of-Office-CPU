module ID_Stage(
    
);


endmodule