module ID_Stage(
    input if_id_stage_reg_t if_id_stage_reg,
    output 
);


endmodule